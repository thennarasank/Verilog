//design
module 2to1_mux
(input i0,i1,s, output y);
assign
assign
endmodule

//test_bench
